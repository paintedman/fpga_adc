
module pll (
	inclk,
	outclk);	

	input		inclk;
	output		outclk;
endmodule
